// nios_qsys.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module nios_qsys (
		input  wire        clk_clk,                                              //                                 clk.clk
		output wire [7:0]  led_pio_export,                                       //                             led_pio.export
		inout  wire        light_i2c_opencores_export_scl_pad_io,                //          light_i2c_opencores_export.scl_pad_io
		inout  wire        light_i2c_opencores_export_sda_pad_io,                //                                    .sda_pad_io
		input  wire        light_int_external_connection_export,                 //       light_int_external_connection.export
		output wire        mm_bridge_for_hps_s0_waitrequest,                     //                mm_bridge_for_hps_s0.waitrequest
		output wire [31:0] mm_bridge_for_hps_s0_readdata,                        //                                    .readdata
		output wire        mm_bridge_for_hps_s0_readdatavalid,                   //                                    .readdatavalid
		input  wire [0:0]  mm_bridge_for_hps_s0_burstcount,                      //                                    .burstcount
		input  wire [31:0] mm_bridge_for_hps_s0_writedata,                       //                                    .writedata
		input  wire [17:0] mm_bridge_for_hps_s0_address,                         //                                    .address
		input  wire        mm_bridge_for_hps_s0_write,                           //                                    .write
		input  wire        mm_bridge_for_hps_s0_read,                            //                                    .read
		input  wire [3:0]  mm_bridge_for_hps_s0_byteenable,                      //                                    .byteenable
		input  wire        mm_bridge_for_hps_s0_debugaccess,                     //                                    .debugaccess
		inout  wire        mpu_i2c_opencores_export_scl_pad_io,                  //            mpu_i2c_opencores_export.scl_pad_io
		inout  wire        mpu_i2c_opencores_export_sda_pad_io,                  //                                    .sda_pad_io
		input  wire        mpu_int_external_connection_export,                   //         mpu_int_external_connection.export
		input  wire        nios2_gen2_cpu_resetrequest_conduit_cpu_resetrequest, // nios2_gen2_cpu_resetrequest_conduit.cpu_resetrequest
		output wire        nios2_gen2_cpu_resetrequest_conduit_cpu_resettaken,   //                                    .cpu_resettaken
		input  wire        reset_reset_n,                                        //                               reset.reset_n
		input  wire        rh_temp_drdy_n_external_connection_export,            //  rh_temp_drdy_n_external_connection.export
		inout  wire        rh_temp_i2c_opencores_export_scl_pad_io,              //        rh_temp_i2c_opencores_export.scl_pad_io
		inout  wire        rh_temp_i2c_opencores_export_sda_pad_io,              //                                    .sda_pad_io
		input  wire        spi_analog_external_MISO,                             //                 spi_analog_external.MISO
		output wire        spi_analog_external_MOSI,                             //                                    .MOSI
		output wire        spi_analog_external_SCLK,                             //                                    .SCLK
		output wire [3:0]  spi_analog_external_SS_n                              //                                    .SS_n
	);

	wire  [31:0] nios2_gen2_data_master_readdata;                                    // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                                 // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                                 // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [18:0] nios2_gen2_data_master_address;                                     // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                                  // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                                        // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_write;                                       // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                                   // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                             // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                          // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [18:0] nios2_gen2_instruction_master_address;                              // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                                 // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         mm_bridge_for_hps_m0_waitrequest;                                   // mm_interconnect_0:mm_bridge_for_hps_m0_waitrequest -> mm_bridge_for_hps:m0_waitrequest
	wire  [31:0] mm_bridge_for_hps_m0_readdata;                                      // mm_interconnect_0:mm_bridge_for_hps_m0_readdata -> mm_bridge_for_hps:m0_readdata
	wire         mm_bridge_for_hps_m0_debugaccess;                                   // mm_bridge_for_hps:m0_debugaccess -> mm_interconnect_0:mm_bridge_for_hps_m0_debugaccess
	wire  [17:0] mm_bridge_for_hps_m0_address;                                       // mm_bridge_for_hps:m0_address -> mm_interconnect_0:mm_bridge_for_hps_m0_address
	wire         mm_bridge_for_hps_m0_read;                                          // mm_bridge_for_hps:m0_read -> mm_interconnect_0:mm_bridge_for_hps_m0_read
	wire   [3:0] mm_bridge_for_hps_m0_byteenable;                                    // mm_bridge_for_hps:m0_byteenable -> mm_interconnect_0:mm_bridge_for_hps_m0_byteenable
	wire         mm_bridge_for_hps_m0_readdatavalid;                                 // mm_interconnect_0:mm_bridge_for_hps_m0_readdatavalid -> mm_bridge_for_hps:m0_readdatavalid
	wire  [31:0] mm_bridge_for_hps_m0_writedata;                                     // mm_bridge_for_hps:m0_writedata -> mm_interconnect_0:mm_bridge_for_hps_m0_writedata
	wire         mm_bridge_for_hps_m0_write;                                         // mm_bridge_for_hps:m0_write -> mm_interconnect_0:mm_bridge_for_hps_m0_write
	wire   [0:0] mm_bridge_for_hps_m0_burstcount;                                    // mm_bridge_for_hps:m0_burstcount -> mm_interconnect_0:mm_bridge_for_hps_m0_burstcount
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;             // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;          // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_chipselect;      // mm_interconnect_0:mpu_i2c_opencores_avalon_slave_0_chipselect -> mpu_i2c_opencores:wb_stb_i
	wire   [7:0] mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_readdata;        // mpu_i2c_opencores:wb_dat_o -> mm_interconnect_0:mpu_i2c_opencores_avalon_slave_0_readdata
	wire         mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_waitrequest;     // mpu_i2c_opencores:wb_ack_o -> mm_interconnect_0:mpu_i2c_opencores_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_address;         // mm_interconnect_0:mpu_i2c_opencores_avalon_slave_0_address -> mpu_i2c_opencores:wb_adr_i
	wire         mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_write;           // mm_interconnect_0:mpu_i2c_opencores_avalon_slave_0_write -> mpu_i2c_opencores:wb_we_i
	wire   [7:0] mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_writedata;       // mm_interconnect_0:mpu_i2c_opencores_avalon_slave_0_writedata -> mpu_i2c_opencores:wb_dat_i
	wire         mm_interconnect_0_light_i2c_opencores_avalon_slave_0_chipselect;    // mm_interconnect_0:light_i2c_opencores_avalon_slave_0_chipselect -> light_i2c_opencores:wb_stb_i
	wire   [7:0] mm_interconnect_0_light_i2c_opencores_avalon_slave_0_readdata;      // light_i2c_opencores:wb_dat_o -> mm_interconnect_0:light_i2c_opencores_avalon_slave_0_readdata
	wire         mm_interconnect_0_light_i2c_opencores_avalon_slave_0_waitrequest;   // light_i2c_opencores:wb_ack_o -> mm_interconnect_0:light_i2c_opencores_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_light_i2c_opencores_avalon_slave_0_address;       // mm_interconnect_0:light_i2c_opencores_avalon_slave_0_address -> light_i2c_opencores:wb_adr_i
	wire         mm_interconnect_0_light_i2c_opencores_avalon_slave_0_write;         // mm_interconnect_0:light_i2c_opencores_avalon_slave_0_write -> light_i2c_opencores:wb_we_i
	wire   [7:0] mm_interconnect_0_light_i2c_opencores_avalon_slave_0_writedata;     // mm_interconnect_0:light_i2c_opencores_avalon_slave_0_writedata -> light_i2c_opencores:wb_dat_i
	wire         mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_chipselect;  // mm_interconnect_0:rh_temp_i2c_opencores_avalon_slave_0_chipselect -> rh_temp_i2c_opencores:wb_stb_i
	wire   [7:0] mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_readdata;    // rh_temp_i2c_opencores:wb_dat_o -> mm_interconnect_0:rh_temp_i2c_opencores_avalon_slave_0_readdata
	wire         mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_waitrequest; // rh_temp_i2c_opencores:wb_ack_o -> mm_interconnect_0:rh_temp_i2c_opencores_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_address;     // mm_interconnect_0:rh_temp_i2c_opencores_avalon_slave_0_address -> rh_temp_i2c_opencores:wb_adr_i
	wire         mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_write;       // mm_interconnect_0:rh_temp_i2c_opencores_avalon_slave_0_write -> rh_temp_i2c_opencores:wb_we_i
	wire   [7:0] mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_writedata;   // mm_interconnect_0:rh_temp_i2c_opencores_avalon_slave_0_writedata -> rh_temp_i2c_opencores:wb_dat_i
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;                // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                 // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;              // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;           // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;           // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;               // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;                  // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;            // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;                 // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;             // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                     // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                       // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_s1_address;                        // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                     // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                          // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                      // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                          // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                              // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                 // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                   // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                               // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_mpu_int_s1_chipselect;                            // mm_interconnect_0:mpu_int_s1_chipselect -> mpu_int:chipselect
	wire  [31:0] mm_interconnect_0_mpu_int_s1_readdata;                              // mpu_int:readdata -> mm_interconnect_0:mpu_int_s1_readdata
	wire   [1:0] mm_interconnect_0_mpu_int_s1_address;                               // mm_interconnect_0:mpu_int_s1_address -> mpu_int:address
	wire         mm_interconnect_0_mpu_int_s1_write;                                 // mm_interconnect_0:mpu_int_s1_write -> mpu_int:write_n
	wire  [31:0] mm_interconnect_0_mpu_int_s1_writedata;                             // mm_interconnect_0:mpu_int_s1_writedata -> mpu_int:writedata
	wire         mm_interconnect_0_light_int_s1_chipselect;                          // mm_interconnect_0:light_int_s1_chipselect -> light_int:chipselect
	wire  [31:0] mm_interconnect_0_light_int_s1_readdata;                            // light_int:readdata -> mm_interconnect_0:light_int_s1_readdata
	wire   [1:0] mm_interconnect_0_light_int_s1_address;                             // mm_interconnect_0:light_int_s1_address -> light_int:address
	wire         mm_interconnect_0_light_int_s1_write;                               // mm_interconnect_0:light_int_s1_write -> light_int:write_n
	wire  [31:0] mm_interconnect_0_light_int_s1_writedata;                           // mm_interconnect_0:light_int_s1_writedata -> light_int:writedata
	wire  [31:0] mm_interconnect_0_rh_temp_drdy_n_s1_readdata;                       // rh_temp_drdy_n:readdata -> mm_interconnect_0:rh_temp_drdy_n_s1_readdata
	wire   [1:0] mm_interconnect_0_rh_temp_drdy_n_s1_address;                        // mm_interconnect_0:rh_temp_drdy_n_s1_address -> rh_temp_drdy_n:address
	wire         mm_interconnect_0_led_pio_s1_chipselect;                            // mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_0_led_pio_s1_readdata;                              // led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_led_pio_s1_address;                               // mm_interconnect_0:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_0_led_pio_s1_write;                                 // mm_interconnect_0:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_0_led_pio_s1_writedata;                             // mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	wire         mm_interconnect_0_shared_memory_s1_chipselect;                      // mm_interconnect_0:shared_memory_s1_chipselect -> shared_memory:chipselect
	wire  [31:0] mm_interconnect_0_shared_memory_s1_readdata;                        // shared_memory:readdata -> mm_interconnect_0:shared_memory_s1_readdata
	wire   [9:0] mm_interconnect_0_shared_memory_s1_address;                         // mm_interconnect_0:shared_memory_s1_address -> shared_memory:address
	wire   [3:0] mm_interconnect_0_shared_memory_s1_byteenable;                      // mm_interconnect_0:shared_memory_s1_byteenable -> shared_memory:byteenable
	wire         mm_interconnect_0_shared_memory_s1_write;                           // mm_interconnect_0:shared_memory_s1_write -> shared_memory:write
	wire  [31:0] mm_interconnect_0_shared_memory_s1_writedata;                       // mm_interconnect_0:shared_memory_s1_writedata -> shared_memory:writedata
	wire         mm_interconnect_0_shared_memory_s1_clken;                           // mm_interconnect_0:shared_memory_s1_clken -> shared_memory:clken
	wire         mm_interconnect_0_spi_analog_spi_control_port_chipselect;           // mm_interconnect_0:spi_analog_spi_control_port_chipselect -> spi_analog:spi_select
	wire  [15:0] mm_interconnect_0_spi_analog_spi_control_port_readdata;             // spi_analog:data_to_cpu -> mm_interconnect_0:spi_analog_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_analog_spi_control_port_address;              // mm_interconnect_0:spi_analog_spi_control_port_address -> spi_analog:mem_addr
	wire         mm_interconnect_0_spi_analog_spi_control_port_read;                 // mm_interconnect_0:spi_analog_spi_control_port_read -> spi_analog:read_n
	wire         mm_interconnect_0_spi_analog_spi_control_port_write;                // mm_interconnect_0:spi_analog_spi_control_port_write -> spi_analog:write_n
	wire  [15:0] mm_interconnect_0_spi_analog_spi_control_port_writedata;            // mm_interconnect_0:spi_analog_spi_control_port_writedata -> spi_analog:data_from_cpu
	wire         mm_interconnect_0_shared_memory_s2_chipselect;                      // mm_interconnect_0:shared_memory_s2_chipselect -> shared_memory:chipselect2
	wire  [31:0] mm_interconnect_0_shared_memory_s2_readdata;                        // shared_memory:readdata2 -> mm_interconnect_0:shared_memory_s2_readdata
	wire   [9:0] mm_interconnect_0_shared_memory_s2_address;                         // mm_interconnect_0:shared_memory_s2_address -> shared_memory:address2
	wire   [3:0] mm_interconnect_0_shared_memory_s2_byteenable;                      // mm_interconnect_0:shared_memory_s2_byteenable -> shared_memory:byteenable2
	wire         mm_interconnect_0_shared_memory_s2_write;                           // mm_interconnect_0:shared_memory_s2_write -> shared_memory:write2
	wire  [31:0] mm_interconnect_0_shared_memory_s2_writedata;                       // mm_interconnect_0:shared_memory_s2_writedata -> shared_memory:writedata2
	wire         mm_interconnect_0_shared_memory_s2_clken;                           // mm_interconnect_0:shared_memory_s2_clken -> shared_memory:clken2
	wire         irq_mapper_receiver0_irq;                                           // mpu_i2c_opencores:wb_inta_o -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                           // light_i2c_opencores:wb_inta_o -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                           // rh_temp_i2c_opencores:wb_inta_o -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                           // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                           // timer:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                           // mpu_int:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                           // light_int:irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                           // spi_analog:irq -> irq_mapper:receiver7_irq
	wire  [31:0] nios2_gen2_irq_irq;                                                 // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [jtag_uart:rst_n, led_pio:reset_n, light_i2c_opencores:wb_rst_i, light_int:reset_n, mm_bridge_for_hps:reset, mm_interconnect_0:mm_bridge_for_hps_reset_reset_bridge_in_reset_reset, mpu_i2c_opencores:wb_rst_i, mpu_int:reset_n, onchip_memory2:reset, rh_temp_drdy_n:reset_n, rh_temp_i2c_opencores:wb_rst_i, rst_translator:in_reset, shared_memory:reset, spi_analog:reset_n, sysid_qsys:reset_n, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                                 // rst_controller:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in, shared_memory:reset_req]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                             // rst_controller_001:reset_req -> [nios2_gen2:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_debug_reset_request_reset;                               // nios2_gen2:debug_reset_request -> rst_controller_001:reset_in1

	nios_qsys_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	nios_qsys_led_pio led_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_export)                           // external_connection.export
	);

	i2c_opencores light_i2c_opencores (
		.wb_clk_i   (clk_clk),                                                          //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                   //      clock_reset.reset
		.scl_pad_io (light_i2c_opencores_export_scl_pad_io),                            //           export.export
		.sda_pad_io (light_i2c_opencores_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver1_irq)                                          // interrupt_sender.irq
	);

	nios_qsys_light_int light_int (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_light_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_light_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_light_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_light_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_light_int_s1_readdata),   //                    .readdata
		.in_port    (light_int_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver6_irq)                   //                 irq.irq
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (18),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_for_hps (
		.clk              (clk_clk),                            //   clk.clk
		.reset            (rst_controller_reset_out_reset),     // reset.reset
		.s0_waitrequest   (mm_bridge_for_hps_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_bridge_for_hps_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_bridge_for_hps_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_bridge_for_hps_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_bridge_for_hps_s0_writedata),     //      .writedata
		.s0_address       (mm_bridge_for_hps_s0_address),       //      .address
		.s0_write         (mm_bridge_for_hps_s0_write),         //      .write
		.s0_read          (mm_bridge_for_hps_s0_read),          //      .read
		.s0_byteenable    (mm_bridge_for_hps_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_bridge_for_hps_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_for_hps_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (mm_bridge_for_hps_m0_readdata),      //      .readdata
		.m0_readdatavalid (mm_bridge_for_hps_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (mm_bridge_for_hps_m0_burstcount),    //      .burstcount
		.m0_writedata     (mm_bridge_for_hps_m0_writedata),     //      .writedata
		.m0_address       (mm_bridge_for_hps_m0_address),       //      .address
		.m0_write         (mm_bridge_for_hps_m0_write),         //      .write
		.m0_read          (mm_bridge_for_hps_m0_read),          //      .read
		.m0_byteenable    (mm_bridge_for_hps_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (mm_bridge_for_hps_m0_debugaccess),   //      .debugaccess
		.s0_response      (),                                   // (terminated)
		.m0_response      (2'b00)                               // (terminated)
	);

	i2c_opencores mpu_i2c_opencores (
		.wb_clk_i   (clk_clk),                                                        //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                 //      clock_reset.reset
		.scl_pad_io (mpu_i2c_opencores_export_scl_pad_io),                            //           export.export
		.sda_pad_io (mpu_i2c_opencores_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver0_irq)                                        // interrupt_sender.irq
	);

	nios_qsys_light_int mpu_int (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_mpu_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mpu_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mpu_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mpu_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mpu_int_s1_readdata),   //                    .readdata
		.in_port    (mpu_int_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                 //                 irq.irq
	);

	nios_qsys_nios2_gen2 nios2_gen2 (
		.clk                                 (clk_clk),                                                  //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       (),                                                         // custom_instruction_master.readra
		.cpu_resetrequest                    (nios2_gen2_cpu_resetrequest_conduit_cpu_resetrequest),     //  cpu_resetrequest_conduit.cpu_resetrequest
		.cpu_resettaken                      (nios2_gen2_cpu_resetrequest_conduit_cpu_resettaken)        //                          .cpu_resettaken
	);

	nios_qsys_onchip_memory2 onchip_memory2 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	nios_qsys_rh_temp_drdy_n rh_temp_drdy_n (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_rh_temp_drdy_n_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_rh_temp_drdy_n_s1_readdata), //                    .readdata
		.in_port  (rh_temp_drdy_n_external_connection_export)     // external_connection.export
	);

	i2c_opencores rh_temp_i2c_opencores (
		.wb_clk_i   (clk_clk),                                                            //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                     //      clock_reset.reset
		.scl_pad_io (rh_temp_i2c_opencores_export_scl_pad_io),                            //           export.export
		.sda_pad_io (rh_temp_i2c_opencores_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver2_irq)                                            // interrupt_sender.irq
	);

	nios_qsys_shared_memory shared_memory (
		.address     (mm_interconnect_0_shared_memory_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_shared_memory_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_shared_memory_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_shared_memory_s1_write),      //       .write
		.readdata    (mm_interconnect_0_shared_memory_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_shared_memory_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_shared_memory_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_shared_memory_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_shared_memory_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_shared_memory_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_shared_memory_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_shared_memory_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_shared_memory_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_shared_memory_s2_byteenable), //       .byteenable
		.clk         (clk_clk),                                       //   clk1.clk
		.reset       (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze      (1'b0)                                           // (terminated)
	);

	nios_qsys_spi_analog spi_analog (
		.clk           (clk_clk),                                                  //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                          //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_analog_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_analog_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_analog_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_analog_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_analog_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_analog_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver7_irq),                                 //              irq.irq
		.MISO          (spi_analog_external_MISO),                                 //         external.export
		.MOSI          (spi_analog_external_MOSI),                                 //                 .export
		.SCLK          (spi_analog_external_SCLK),                                 //                 .export
		.SS_n          (spi_analog_external_SS_n)                                  //                 .export
	);

	nios_qsys_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	nios_qsys_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)               //   irq.irq
	);

	nios_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                      (clk_clk),                                                             //                                    clk_50_clk.clk
		.mm_bridge_for_hps_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                      // mm_bridge_for_hps_reset_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                                  //        nios2_gen2_reset_reset_bridge_in_reset.reset
		.mm_bridge_for_hps_m0_address                        (mm_bridge_for_hps_m0_address),                                        //                          mm_bridge_for_hps_m0.address
		.mm_bridge_for_hps_m0_waitrequest                    (mm_bridge_for_hps_m0_waitrequest),                                    //                                              .waitrequest
		.mm_bridge_for_hps_m0_burstcount                     (mm_bridge_for_hps_m0_burstcount),                                     //                                              .burstcount
		.mm_bridge_for_hps_m0_byteenable                     (mm_bridge_for_hps_m0_byteenable),                                     //                                              .byteenable
		.mm_bridge_for_hps_m0_read                           (mm_bridge_for_hps_m0_read),                                           //                                              .read
		.mm_bridge_for_hps_m0_readdata                       (mm_bridge_for_hps_m0_readdata),                                       //                                              .readdata
		.mm_bridge_for_hps_m0_readdatavalid                  (mm_bridge_for_hps_m0_readdatavalid),                                  //                                              .readdatavalid
		.mm_bridge_for_hps_m0_write                          (mm_bridge_for_hps_m0_write),                                          //                                              .write
		.mm_bridge_for_hps_m0_writedata                      (mm_bridge_for_hps_m0_writedata),                                      //                                              .writedata
		.mm_bridge_for_hps_m0_debugaccess                    (mm_bridge_for_hps_m0_debugaccess),                                    //                                              .debugaccess
		.nios2_gen2_data_master_address                      (nios2_gen2_data_master_address),                                      //                        nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                  (nios2_gen2_data_master_waitrequest),                                  //                                              .waitrequest
		.nios2_gen2_data_master_byteenable                   (nios2_gen2_data_master_byteenable),                                   //                                              .byteenable
		.nios2_gen2_data_master_read                         (nios2_gen2_data_master_read),                                         //                                              .read
		.nios2_gen2_data_master_readdata                     (nios2_gen2_data_master_readdata),                                     //                                              .readdata
		.nios2_gen2_data_master_write                        (nios2_gen2_data_master_write),                                        //                                              .write
		.nios2_gen2_data_master_writedata                    (nios2_gen2_data_master_writedata),                                    //                                              .writedata
		.nios2_gen2_data_master_debugaccess                  (nios2_gen2_data_master_debugaccess),                                  //                                              .debugaccess
		.nios2_gen2_instruction_master_address               (nios2_gen2_instruction_master_address),                               //                 nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest           (nios2_gen2_instruction_master_waitrequest),                           //                                              .waitrequest
		.nios2_gen2_instruction_master_read                  (nios2_gen2_instruction_master_read),                                  //                                              .read
		.nios2_gen2_instruction_master_readdata              (nios2_gen2_instruction_master_readdata),                              //                                              .readdata
		.jtag_uart_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),               //                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                 //                                              .write
		.jtag_uart_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                  //                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),              //                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),             //                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),           //                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),            //                                              .chipselect
		.led_pio_s1_address                                  (mm_interconnect_0_led_pio_s1_address),                                //                                    led_pio_s1.address
		.led_pio_s1_write                                    (mm_interconnect_0_led_pio_s1_write),                                  //                                              .write
		.led_pio_s1_readdata                                 (mm_interconnect_0_led_pio_s1_readdata),                               //                                              .readdata
		.led_pio_s1_writedata                                (mm_interconnect_0_led_pio_s1_writedata),                              //                                              .writedata
		.led_pio_s1_chipselect                               (mm_interconnect_0_led_pio_s1_chipselect),                             //                                              .chipselect
		.light_i2c_opencores_avalon_slave_0_address          (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_address),        //            light_i2c_opencores_avalon_slave_0.address
		.light_i2c_opencores_avalon_slave_0_write            (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_write),          //                                              .write
		.light_i2c_opencores_avalon_slave_0_readdata         (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_readdata),       //                                              .readdata
		.light_i2c_opencores_avalon_slave_0_writedata        (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_writedata),      //                                              .writedata
		.light_i2c_opencores_avalon_slave_0_waitrequest      (~mm_interconnect_0_light_i2c_opencores_avalon_slave_0_waitrequest),   //                                              .waitrequest
		.light_i2c_opencores_avalon_slave_0_chipselect       (mm_interconnect_0_light_i2c_opencores_avalon_slave_0_chipselect),     //                                              .chipselect
		.light_int_s1_address                                (mm_interconnect_0_light_int_s1_address),                              //                                  light_int_s1.address
		.light_int_s1_write                                  (mm_interconnect_0_light_int_s1_write),                                //                                              .write
		.light_int_s1_readdata                               (mm_interconnect_0_light_int_s1_readdata),                             //                                              .readdata
		.light_int_s1_writedata                              (mm_interconnect_0_light_int_s1_writedata),                            //                                              .writedata
		.light_int_s1_chipselect                             (mm_interconnect_0_light_int_s1_chipselect),                           //                                              .chipselect
		.mpu_i2c_opencores_avalon_slave_0_address            (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_address),          //              mpu_i2c_opencores_avalon_slave_0.address
		.mpu_i2c_opencores_avalon_slave_0_write              (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_write),            //                                              .write
		.mpu_i2c_opencores_avalon_slave_0_readdata           (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_readdata),         //                                              .readdata
		.mpu_i2c_opencores_avalon_slave_0_writedata          (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_writedata),        //                                              .writedata
		.mpu_i2c_opencores_avalon_slave_0_waitrequest        (~mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_waitrequest),     //                                              .waitrequest
		.mpu_i2c_opencores_avalon_slave_0_chipselect         (mm_interconnect_0_mpu_i2c_opencores_avalon_slave_0_chipselect),       //                                              .chipselect
		.mpu_int_s1_address                                  (mm_interconnect_0_mpu_int_s1_address),                                //                                    mpu_int_s1.address
		.mpu_int_s1_write                                    (mm_interconnect_0_mpu_int_s1_write),                                  //                                              .write
		.mpu_int_s1_readdata                                 (mm_interconnect_0_mpu_int_s1_readdata),                               //                                              .readdata
		.mpu_int_s1_writedata                                (mm_interconnect_0_mpu_int_s1_writedata),                              //                                              .writedata
		.mpu_int_s1_chipselect                               (mm_interconnect_0_mpu_int_s1_chipselect),                             //                                              .chipselect
		.nios2_gen2_debug_mem_slave_address                  (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),                //                    nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                    (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),                  //                                              .write
		.nios2_gen2_debug_mem_slave_read                     (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),                   //                                              .read
		.nios2_gen2_debug_mem_slave_readdata                 (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),               //                                              .readdata
		.nios2_gen2_debug_mem_slave_writedata                (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),              //                                              .writedata
		.nios2_gen2_debug_mem_slave_byteenable               (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),             //                                              .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest              (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),            //                                              .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess              (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),            //                                              .debugaccess
		.onchip_memory2_s1_address                           (mm_interconnect_0_onchip_memory2_s1_address),                         //                             onchip_memory2_s1.address
		.onchip_memory2_s1_write                             (mm_interconnect_0_onchip_memory2_s1_write),                           //                                              .write
		.onchip_memory2_s1_readdata                          (mm_interconnect_0_onchip_memory2_s1_readdata),                        //                                              .readdata
		.onchip_memory2_s1_writedata                         (mm_interconnect_0_onchip_memory2_s1_writedata),                       //                                              .writedata
		.onchip_memory2_s1_byteenable                        (mm_interconnect_0_onchip_memory2_s1_byteenable),                      //                                              .byteenable
		.onchip_memory2_s1_chipselect                        (mm_interconnect_0_onchip_memory2_s1_chipselect),                      //                                              .chipselect
		.onchip_memory2_s1_clken                             (mm_interconnect_0_onchip_memory2_s1_clken),                           //                                              .clken
		.rh_temp_drdy_n_s1_address                           (mm_interconnect_0_rh_temp_drdy_n_s1_address),                         //                             rh_temp_drdy_n_s1.address
		.rh_temp_drdy_n_s1_readdata                          (mm_interconnect_0_rh_temp_drdy_n_s1_readdata),                        //                                              .readdata
		.rh_temp_i2c_opencores_avalon_slave_0_address        (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_address),      //          rh_temp_i2c_opencores_avalon_slave_0.address
		.rh_temp_i2c_opencores_avalon_slave_0_write          (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_write),        //                                              .write
		.rh_temp_i2c_opencores_avalon_slave_0_readdata       (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_readdata),     //                                              .readdata
		.rh_temp_i2c_opencores_avalon_slave_0_writedata      (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_writedata),    //                                              .writedata
		.rh_temp_i2c_opencores_avalon_slave_0_waitrequest    (~mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_waitrequest), //                                              .waitrequest
		.rh_temp_i2c_opencores_avalon_slave_0_chipselect     (mm_interconnect_0_rh_temp_i2c_opencores_avalon_slave_0_chipselect),   //                                              .chipselect
		.shared_memory_s1_address                            (mm_interconnect_0_shared_memory_s1_address),                          //                              shared_memory_s1.address
		.shared_memory_s1_write                              (mm_interconnect_0_shared_memory_s1_write),                            //                                              .write
		.shared_memory_s1_readdata                           (mm_interconnect_0_shared_memory_s1_readdata),                         //                                              .readdata
		.shared_memory_s1_writedata                          (mm_interconnect_0_shared_memory_s1_writedata),                        //                                              .writedata
		.shared_memory_s1_byteenable                         (mm_interconnect_0_shared_memory_s1_byteenable),                       //                                              .byteenable
		.shared_memory_s1_chipselect                         (mm_interconnect_0_shared_memory_s1_chipselect),                       //                                              .chipselect
		.shared_memory_s1_clken                              (mm_interconnect_0_shared_memory_s1_clken),                            //                                              .clken
		.shared_memory_s2_address                            (mm_interconnect_0_shared_memory_s2_address),                          //                              shared_memory_s2.address
		.shared_memory_s2_write                              (mm_interconnect_0_shared_memory_s2_write),                            //                                              .write
		.shared_memory_s2_readdata                           (mm_interconnect_0_shared_memory_s2_readdata),                         //                                              .readdata
		.shared_memory_s2_writedata                          (mm_interconnect_0_shared_memory_s2_writedata),                        //                                              .writedata
		.shared_memory_s2_byteenable                         (mm_interconnect_0_shared_memory_s2_byteenable),                       //                                              .byteenable
		.shared_memory_s2_chipselect                         (mm_interconnect_0_shared_memory_s2_chipselect),                       //                                              .chipselect
		.shared_memory_s2_clken                              (mm_interconnect_0_shared_memory_s2_clken),                            //                                              .clken
		.spi_analog_spi_control_port_address                 (mm_interconnect_0_spi_analog_spi_control_port_address),               //                   spi_analog_spi_control_port.address
		.spi_analog_spi_control_port_write                   (mm_interconnect_0_spi_analog_spi_control_port_write),                 //                                              .write
		.spi_analog_spi_control_port_read                    (mm_interconnect_0_spi_analog_spi_control_port_read),                  //                                              .read
		.spi_analog_spi_control_port_readdata                (mm_interconnect_0_spi_analog_spi_control_port_readdata),              //                                              .readdata
		.spi_analog_spi_control_port_writedata               (mm_interconnect_0_spi_analog_spi_control_port_writedata),             //                                              .writedata
		.spi_analog_spi_control_port_chipselect              (mm_interconnect_0_spi_analog_spi_control_port_chipselect),            //                                              .chipselect
		.sysid_qsys_control_slave_address                    (mm_interconnect_0_sysid_qsys_control_slave_address),                  //                      sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                   (mm_interconnect_0_sysid_qsys_control_slave_readdata),                 //                                              .readdata
		.timer_s1_address                                    (mm_interconnect_0_timer_s1_address),                                  //                                      timer_s1.address
		.timer_s1_write                                      (mm_interconnect_0_timer_s1_write),                                    //                                              .write
		.timer_s1_readdata                                   (mm_interconnect_0_timer_s1_readdata),                                 //                                              .readdata
		.timer_s1_writedata                                  (mm_interconnect_0_timer_s1_writedata),                                //                                              .writedata
		.timer_s1_chipselect                                 (mm_interconnect_0_timer_s1_chipselect)                                //                                              .chipselect
	);

	nios_qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),           // receiver7.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
